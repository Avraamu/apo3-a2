library IEEE;
use IEEE.std_logic_1164.ALL;

entity time is
end time;


