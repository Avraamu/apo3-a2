configuration lanespd_fsm_behaviour_cfg of lanespd_fsm is
   for behaviour
   end for;
end lanespd_fsm_behaviour_cfg;


