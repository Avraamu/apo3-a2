library IEEE;
use IEEE.std_logic_1164.ALL;

entity score is
end score;


