configuration bulletspd_fsm_synthesised_cfg of bulletspd_fsm is
   for synthesised
   end for;
end bulletspd_fsm_synthesised_cfg;


