configuration timebase_synthesised_cfg of timebase is
   for synthesised
   end for;
end timebase_synthesised_cfg;


