configuration bulletspd_fsm_behaviour_cfg of bulletspd_fsm is
   for behaviour
   end for;
end bulletspd_fsm_behaviour_cfg;


