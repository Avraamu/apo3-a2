configuration timebase_behaviour_cfg of timebase is
   for behaviour
   end for;
end timebase_behaviour_cfg;


