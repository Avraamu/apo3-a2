library IEEE;
use IEEE.std_logic_1164.ALL;

entity tb is
end tb;


