library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of inputbuffer is
begin
end behaviour;


