library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of graphics is
begin
end behaviour;


