library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of controller is
begin
end behaviour;





