library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of player is
begin
end behaviour;


