library IEEE;
use IEEE.std_logic_1164.ALL;

entity bulletspd_fsm is
   port(bulletspd  :in    std_logic;
        bulletspd_p:out   std_logic;
        res      :in    std_logic;
        clk        :in    std_logic);
end bulletspd_fsm;





