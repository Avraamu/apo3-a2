library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of collision is
begin
end behaviour;


