configuration lanespd_fsm_synthesised_cfg of lanespd_fsm is
   for synthesised
   end for;
end lanespd_fsm_synthesised_cfg;


