library IEEE;
use IEEE.std_logic_1164.ALL;

entity rng is
end rng;


